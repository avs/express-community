      module libSTM<build_dir="xp_comm_proj/stm/src/lib",process="express",c_src_files="fgetPlainCoord.c fgetSurface.c fgetchem_3d.c fgetcoord.c fgetcube.c fgetdcar.c fgetdmol_xyz.c fgetespcoord.c fgetgamess.c fgetmm3.c fgetmol.c fgetmol2.c fgetmopac.c fgetpdb.c fgetCgamess.c makeatomamin.c makeatomtype.c makeatomtype_prot.c makebonds.c makemainchain.c",c_hdr_files="geomcoord.h">;
